// nios_cpu.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module nios_cpu (
		input  wire        clk_clk,          //       clk.clk
		output wire [7:0]  led_green_export, // led_green.export
		output wire [17:0] led_red_export,   //   led_red.export
		input  wire [3:0]  push_btns_export, // push_btns.export
		input  wire        reset_reset_n,    //     reset.reset_n
		input  wire [17:0] switches_export   //  switches.export
	);

	wire  [31:0] nios_cpu_data_master_readdata;                             // mm_interconnect_0:nios_cpu_data_master_readdata -> nios_cpu:d_readdata
	wire         nios_cpu_data_master_waitrequest;                          // mm_interconnect_0:nios_cpu_data_master_waitrequest -> nios_cpu:d_waitrequest
	wire         nios_cpu_data_master_debugaccess;                          // nios_cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios_cpu_data_master_debugaccess
	wire  [19:0] nios_cpu_data_master_address;                              // nios_cpu:d_address -> mm_interconnect_0:nios_cpu_data_master_address
	wire   [3:0] nios_cpu_data_master_byteenable;                           // nios_cpu:d_byteenable -> mm_interconnect_0:nios_cpu_data_master_byteenable
	wire         nios_cpu_data_master_read;                                 // nios_cpu:d_read -> mm_interconnect_0:nios_cpu_data_master_read
	wire         nios_cpu_data_master_readdatavalid;                        // mm_interconnect_0:nios_cpu_data_master_readdatavalid -> nios_cpu:d_readdatavalid
	wire         nios_cpu_data_master_write;                                // nios_cpu:d_write -> mm_interconnect_0:nios_cpu_data_master_write
	wire  [31:0] nios_cpu_data_master_writedata;                            // nios_cpu:d_writedata -> mm_interconnect_0:nios_cpu_data_master_writedata
	wire  [31:0] nios_cpu_instruction_master_readdata;                      // mm_interconnect_0:nios_cpu_instruction_master_readdata -> nios_cpu:i_readdata
	wire         nios_cpu_instruction_master_waitrequest;                   // mm_interconnect_0:nios_cpu_instruction_master_waitrequest -> nios_cpu:i_waitrequest
	wire  [19:0] nios_cpu_instruction_master_address;                       // nios_cpu:i_address -> mm_interconnect_0:nios_cpu_instruction_master_address
	wire         nios_cpu_instruction_master_read;                          // nios_cpu:i_read -> mm_interconnect_0:nios_cpu_instruction_master_read
	wire         nios_cpu_instruction_master_readdatavalid;                 // mm_interconnect_0:nios_cpu_instruction_master_readdatavalid -> nios_cpu:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;     // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;      // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios_cpu_debug_mem_slave_readdata;       // nios_cpu:debug_mem_slave_readdata -> mm_interconnect_0:nios_cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios_cpu_debug_mem_slave_waitrequest;    // nios_cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:nios_cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios_cpu_debug_mem_slave_debugaccess;    // mm_interconnect_0:nios_cpu_debug_mem_slave_debugaccess -> nios_cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios_cpu_debug_mem_slave_address;        // mm_interconnect_0:nios_cpu_debug_mem_slave_address -> nios_cpu:debug_mem_slave_address
	wire         mm_interconnect_0_nios_cpu_debug_mem_slave_read;           // mm_interconnect_0:nios_cpu_debug_mem_slave_read -> nios_cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios_cpu_debug_mem_slave_byteenable;     // mm_interconnect_0:nios_cpu_debug_mem_slave_byteenable -> nios_cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios_cpu_debug_mem_slave_write;          // mm_interconnect_0:nios_cpu_debug_mem_slave_write -> nios_cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios_cpu_debug_mem_slave_writedata;      // mm_interconnect_0:nios_cpu_debug_mem_slave_writedata -> nios_cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_led_green_s1_chipselect;                 // mm_interconnect_0:led_green_s1_chipselect -> led_green:chipselect
	wire  [31:0] mm_interconnect_0_led_green_s1_readdata;                   // led_green:readdata -> mm_interconnect_0:led_green_s1_readdata
	wire   [1:0] mm_interconnect_0_led_green_s1_address;                    // mm_interconnect_0:led_green_s1_address -> led_green:address
	wire         mm_interconnect_0_led_green_s1_write;                      // mm_interconnect_0:led_green_s1_write -> led_green:write_n
	wire  [31:0] mm_interconnect_0_led_green_s1_writedata;                  // mm_interconnect_0:led_green_s1_writedata -> led_green:writedata
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;             // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;               // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [15:0] mm_interconnect_0_onchip_memory_s1_address;                // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;             // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                  // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;              // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                  // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_led_red_s1_chipselect;                   // mm_interconnect_0:led_red_s1_chipselect -> led_red:chipselect
	wire  [31:0] mm_interconnect_0_led_red_s1_readdata;                     // led_red:readdata -> mm_interconnect_0:led_red_s1_readdata
	wire   [1:0] mm_interconnect_0_led_red_s1_address;                      // mm_interconnect_0:led_red_s1_address -> led_red:address
	wire         mm_interconnect_0_led_red_s1_write;                        // mm_interconnect_0:led_red_s1_write -> led_red:write_n
	wire  [31:0] mm_interconnect_0_led_red_s1_writedata;                    // mm_interconnect_0:led_red_s1_writedata -> led_red:writedata
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;                    // switches:readdata -> mm_interconnect_0:switches_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_s1_address;                     // mm_interconnect_0:switches_s1_address -> switches:address
	wire         mm_interconnect_0_push_btns_s1_chipselect;                 // mm_interconnect_0:push_btns_s1_chipselect -> push_btns:chipselect
	wire  [31:0] mm_interconnect_0_push_btns_s1_readdata;                   // push_btns:readdata -> mm_interconnect_0:push_btns_s1_readdata
	wire   [1:0] mm_interconnect_0_push_btns_s1_address;                    // mm_interconnect_0:push_btns_s1_address -> push_btns:address
	wire         mm_interconnect_0_push_btns_s1_write;                      // mm_interconnect_0:push_btns_s1_write -> push_btns:write_n
	wire  [31:0] mm_interconnect_0_push_btns_s1_writedata;                  // mm_interconnect_0:push_btns_s1_writedata -> push_btns:writedata
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // push_btns:irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios_cpu_irq_irq;                                          // irq_mapper:sender_irq -> nios_cpu:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [irq_mapper:reset, jtag_uart:rst_n, led_green:reset_n, led_red:reset_n, mm_interconnect_0:nios_cpu_reset_reset_bridge_in_reset_reset, nios_cpu:reset_n, onchip_memory:reset, push_btns:reset_n, rst_translator:in_reset, switches:reset_n, sysid_qsys_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [nios_cpu:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	wire         nios_cpu_debug_reset_request_reset;                        // nios_cpu:debug_reset_request -> rst_controller:reset_in1

	nios_cpu_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	nios_cpu_led_green led_green (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_led_green_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_green_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_green_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_green_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_green_s1_readdata),   //                    .readdata
		.out_port   (led_green_export)                           // external_connection.export
	);

	nios_cpu_led_red led_red (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_led_red_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_red_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_red_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_red_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_red_s1_readdata),   //                    .readdata
		.out_port   (led_red_export)                           // external_connection.export
	);

	nios_cpu_nios_cpu nios_cpu (
		.clk                                 (clk_clk),                                                //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios_cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios_cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios_cpu_data_master_read),                              //                          .read
		.d_readdata                          (nios_cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios_cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios_cpu_data_master_write),                             //                          .write
		.d_writedata                         (nios_cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios_cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios_cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios_cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios_cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (nios_cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios_cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios_cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios_cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios_cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                        // custom_instruction_master.readra
	);

	nios_cpu_onchip_memory onchip_memory (
		.clk        (clk_clk),                                       //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),            //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	nios_cpu_push_btns push_btns (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_push_btns_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_push_btns_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_push_btns_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_push_btns_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_push_btns_s1_readdata),   //                    .readdata
		.in_port    (push_btns_export),                          // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                   //                 irq.irq
	);

	nios_cpu_switches switches (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switches_s1_readdata), //                    .readdata
		.in_port  (switches_export)                         // external_connection.export
	);

	nios_cpu_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	nios_cpu_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                             (clk_clk),                                                   //                           clk_50_clk.clk
		.nios_cpu_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // nios_cpu_reset_reset_bridge_in_reset.reset
		.nios_cpu_data_master_address               (nios_cpu_data_master_address),                              //                 nios_cpu_data_master.address
		.nios_cpu_data_master_waitrequest           (nios_cpu_data_master_waitrequest),                          //                                     .waitrequest
		.nios_cpu_data_master_byteenable            (nios_cpu_data_master_byteenable),                           //                                     .byteenable
		.nios_cpu_data_master_read                  (nios_cpu_data_master_read),                                 //                                     .read
		.nios_cpu_data_master_readdata              (nios_cpu_data_master_readdata),                             //                                     .readdata
		.nios_cpu_data_master_readdatavalid         (nios_cpu_data_master_readdatavalid),                        //                                     .readdatavalid
		.nios_cpu_data_master_write                 (nios_cpu_data_master_write),                                //                                     .write
		.nios_cpu_data_master_writedata             (nios_cpu_data_master_writedata),                            //                                     .writedata
		.nios_cpu_data_master_debugaccess           (nios_cpu_data_master_debugaccess),                          //                                     .debugaccess
		.nios_cpu_instruction_master_address        (nios_cpu_instruction_master_address),                       //          nios_cpu_instruction_master.address
		.nios_cpu_instruction_master_waitrequest    (nios_cpu_instruction_master_waitrequest),                   //                                     .waitrequest
		.nios_cpu_instruction_master_read           (nios_cpu_instruction_master_read),                          //                                     .read
		.nios_cpu_instruction_master_readdata       (nios_cpu_instruction_master_readdata),                      //                                     .readdata
		.nios_cpu_instruction_master_readdatavalid  (nios_cpu_instruction_master_readdatavalid),                 //                                     .readdatavalid
		.jtag_uart_avalon_jtag_slave_address        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //          jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                     .write
		.jtag_uart_avalon_jtag_slave_read           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                     .read
		.jtag_uart_avalon_jtag_slave_readdata       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                     .readdata
		.jtag_uart_avalon_jtag_slave_writedata      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                     .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                     .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                     .chipselect
		.led_green_s1_address                       (mm_interconnect_0_led_green_s1_address),                    //                         led_green_s1.address
		.led_green_s1_write                         (mm_interconnect_0_led_green_s1_write),                      //                                     .write
		.led_green_s1_readdata                      (mm_interconnect_0_led_green_s1_readdata),                   //                                     .readdata
		.led_green_s1_writedata                     (mm_interconnect_0_led_green_s1_writedata),                  //                                     .writedata
		.led_green_s1_chipselect                    (mm_interconnect_0_led_green_s1_chipselect),                 //                                     .chipselect
		.led_red_s1_address                         (mm_interconnect_0_led_red_s1_address),                      //                           led_red_s1.address
		.led_red_s1_write                           (mm_interconnect_0_led_red_s1_write),                        //                                     .write
		.led_red_s1_readdata                        (mm_interconnect_0_led_red_s1_readdata),                     //                                     .readdata
		.led_red_s1_writedata                       (mm_interconnect_0_led_red_s1_writedata),                    //                                     .writedata
		.led_red_s1_chipselect                      (mm_interconnect_0_led_red_s1_chipselect),                   //                                     .chipselect
		.nios_cpu_debug_mem_slave_address           (mm_interconnect_0_nios_cpu_debug_mem_slave_address),        //             nios_cpu_debug_mem_slave.address
		.nios_cpu_debug_mem_slave_write             (mm_interconnect_0_nios_cpu_debug_mem_slave_write),          //                                     .write
		.nios_cpu_debug_mem_slave_read              (mm_interconnect_0_nios_cpu_debug_mem_slave_read),           //                                     .read
		.nios_cpu_debug_mem_slave_readdata          (mm_interconnect_0_nios_cpu_debug_mem_slave_readdata),       //                                     .readdata
		.nios_cpu_debug_mem_slave_writedata         (mm_interconnect_0_nios_cpu_debug_mem_slave_writedata),      //                                     .writedata
		.nios_cpu_debug_mem_slave_byteenable        (mm_interconnect_0_nios_cpu_debug_mem_slave_byteenable),     //                                     .byteenable
		.nios_cpu_debug_mem_slave_waitrequest       (mm_interconnect_0_nios_cpu_debug_mem_slave_waitrequest),    //                                     .waitrequest
		.nios_cpu_debug_mem_slave_debugaccess       (mm_interconnect_0_nios_cpu_debug_mem_slave_debugaccess),    //                                     .debugaccess
		.onchip_memory_s1_address                   (mm_interconnect_0_onchip_memory_s1_address),                //                     onchip_memory_s1.address
		.onchip_memory_s1_write                     (mm_interconnect_0_onchip_memory_s1_write),                  //                                     .write
		.onchip_memory_s1_readdata                  (mm_interconnect_0_onchip_memory_s1_readdata),               //                                     .readdata
		.onchip_memory_s1_writedata                 (mm_interconnect_0_onchip_memory_s1_writedata),              //                                     .writedata
		.onchip_memory_s1_byteenable                (mm_interconnect_0_onchip_memory_s1_byteenable),             //                                     .byteenable
		.onchip_memory_s1_chipselect                (mm_interconnect_0_onchip_memory_s1_chipselect),             //                                     .chipselect
		.onchip_memory_s1_clken                     (mm_interconnect_0_onchip_memory_s1_clken),                  //                                     .clken
		.push_btns_s1_address                       (mm_interconnect_0_push_btns_s1_address),                    //                         push_btns_s1.address
		.push_btns_s1_write                         (mm_interconnect_0_push_btns_s1_write),                      //                                     .write
		.push_btns_s1_readdata                      (mm_interconnect_0_push_btns_s1_readdata),                   //                                     .readdata
		.push_btns_s1_writedata                     (mm_interconnect_0_push_btns_s1_writedata),                  //                                     .writedata
		.push_btns_s1_chipselect                    (mm_interconnect_0_push_btns_s1_chipselect),                 //                                     .chipselect
		.switches_s1_address                        (mm_interconnect_0_switches_s1_address),                     //                          switches_s1.address
		.switches_s1_readdata                       (mm_interconnect_0_switches_s1_readdata),                    //                                     .readdata
		.sysid_qsys_0_control_slave_address         (mm_interconnect_0_sysid_qsys_0_control_slave_address),      //           sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata        (mm_interconnect_0_sysid_qsys_0_control_slave_readdata)      //                                     .readdata
	);

	nios_cpu_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios_cpu_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios_cpu_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
